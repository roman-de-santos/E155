module top_tb();